module CU_logic #(parameter states=40) (


    output logic RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,
    PCINC,
    COUNTER_LD,COUNTER_INC,COUNTER_CLR,

    output logic [2:0] ALUSEL,

    output logic [3:0] SYSTEMBUSSEL,

    input logic [states-1:0] CPU_state

);

// must also input NZCV flags
// needed to choose whether to execute the conditional branch instructions or not!


// logic derived in "instructions.txt"

// counter mapping is as follows (40 states - * indicates start state of routine)
// fetch1   : 0
// fetch2   : 1
// fetch3   : 2
// nop1     : 3*
// mov1     : 4*
// ALTmov1  : 5*
// ALTmov2  : 6
// ldr1     : 7*
// ldr2     : 8
// ALTldr1  : 9*
// ALTldr2  : 10
// ALTldr3  : 11
// ALTldr4  : 12
// str1     : 13*
// str2     : 14
// str3     : 15
// str4     : 16
// ALTstr1  : 17*
// ALTstr2  : 18
// ALTstr3  : 19
// ALTstr4  : 20
// cmp1     : 21*
// b1       : 22*
// bgt1     : 23*
// blt1     : 24*
// beq1     : 25*
// add1     : 26*
// add2     : 27
// sub1     : 28*
// sub2     : 29
// mul1     : 30*
// mul2     : 31
// lsr1     : 32*
// lsr2     : 33
// and1     : 34*
// and2     : 35
// or1      : 36*
// or2      : 37
// mvn1     : 38*
// mvn2     : 39


// SYSTEMBUSSEL = 0 : PC
// SYSTEMBUSSEL = 1 : DR
// SYSTEMBUSSEL = 2 : AR
// SYSTEMBUSSEL = 3 : AC
// SYSTEMBUSSEL = 4 : MEM
// SYSTEMBUSSEL = 5 : TR
// SYSTEMBUSSEL = 6 : rop1
// SYSTEMBUSSEL = 7 : rop2
// SYSTEMBUSSEL = 8 : GPR1



always_comb begin

    case(CPU_state)

    40'd2**0 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**1 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**2 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**3 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**4 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**5 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**6 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**7 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**8 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**9 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**10 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**11 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**12 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**13 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**14 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**15 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**16 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**17 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**18 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**19 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**20 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**21 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**22 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**23 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**24 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**25 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**26 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**27 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**28 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**29 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**30 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**31 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**32 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**33 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**34 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**35 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**36 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**37 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**38 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    40'd2**39 : begin
        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;
    end

    default : begin

        {RSELLOAD,ROP1LOAD,ROP2LOAD,TRLOAD,ARLOAD,PCLOAD,DRLOAD,ACLOAD,IRLOAD,GPRLOAD,MEMLOAD,PCINC,COUNTER_LD,COUNTER_INC,COUNTER_CLR} = 'd0;
        ALUSEL = 'd0;
        SYSTEMBUSSEL = 'd0;

    end

    endcase

end











endmodule